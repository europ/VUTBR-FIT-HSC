
//------> C:/PROGRA~1/MENTOR~1/CATAPU~1.0C/Mgc_home/pkgs/siflibs/mgc_in_wire_en_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


`ifdef mgc_in_wire_en_v1
`else
`define mgc_in_wire_en_v1
module mgc_in_wire_en_v1 (ld, d, lz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output [width-1:0] d;
  output             lz;
  input  [width-1:0] z;

  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;

endmodule
`endif


//------> C:/PROGRA~1/MENTOR~1/CATAPU~1.0C/Mgc_home/pkgs/siflibs/mgc_in_wire_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


`ifdef mgc_in_wire_v1
`else
`define mgc_in_wire_v1
module mgc_in_wire_v1 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] d;
  input  [width-1:0] z;

  wire   [width-1:0] d;

  assign d = z;

endmodule
`endif


//------> C:/PROGRA~1/MENTOR~1/CATAPU~1.0C/Mgc_home/pkgs/siflibs/mgc_out_stdreg_en_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


`ifdef mgc_out_stdreg_en_v1
`else
`define mgc_out_stdreg_en_v1
module mgc_out_stdreg_en_v1 (ld, d, lz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  input  [width-1:0] d;
  output             lz;
  output [width-1:0] z;

  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;

endmodule
`endif



//------> C:/PROGRA~1/MENTOR~1/CATAPU~1.0C/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Block 1R1W Read Before Write RAM with common clock
`ifdef BLOCK_1R1W_RBW
`else
`define BLOCK_1R1W_RBW
module BLOCK_1R1W_RBW
#(
parameter data_width = 8,
parameter addr_width = 7,
parameter depth = 128
)(
	radr, wadr, d, we, re, clk, q
);

	input [addr_width-1:0] radr;
	input [addr_width-1:0] wadr;
	input [data_width-1:0] d;
	input we;
	input re;
	input clk;
	output[data_width-1:0] q;

	reg [data_width-1:0] q;

	(* ram_style = "block" *)
	reg [data_width-1:0] mem [depth-1:0];// synthesis syn_ramstyle="block_ram"
	//pragma attribute mem block_ram true
		
	always @(posedge clk) begin
		if (we) begin
			mem[wadr] <= d; // Write port
		end
		if (re) begin
			q <= mem[radr] ; // read port
		end
	end

endmodule
`endif

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0c/745553 Production Release
//  HLS Date:       Wed Oct 11 16:38:17 PDT 2017
// 
//  Generated by:   Fitkit@DESKTOP-NJUNEBJ
//  Generated date: Sat Dec 15 16:31:58 2018
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_3_10_640_7_gen
// ------------------------------------------------------------------


`ifdef Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_3_10_640_7_gen
`else
`define Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_3_10_640_7_gen
module Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_3_10_640_7_gen (
  we, d, wadr, re, q, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d
);
  output we;
  output [2:0] d;
  output [9:0] wadr;
  output re;
  input [2:0] q;
  output [9:0] radr;
  input [9:0] radr_d;
  input [9:0] wadr_d;
  input [2:0] d_d;
  input we_d;
  input re_d;
  output [2:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (we_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule
`endif

// ------------------------------------------------------------------
//  Design Unit:    Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_32_9_512_4_gen
// ------------------------------------------------------------------


`ifdef Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_32_9_512_4_gen
`else
`define Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_32_9_512_4_gen
module Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_32_9_512_4_gen (
  we, d, q, adr, adr_d, d_d, we_d, q_d, ram_rw_A_internal_RMASK_B_d
);
  output we;
  output [31:0] d;
  input [31:0] q;
  output [8:0] adr;
  input [8:0] adr_d;
  input [31:0] d_d;
  input we_d;
  output [31:0] q_d;
  input ram_rw_A_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (we_d);
  assign d = (d_d);
  assign q_d = q;
  assign adr = (adr_d);
endmodule
`endif

// ------------------------------------------------------------------
//  Design Unit:    filter_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


`ifdef filter_core_core_fsm
`else
`define filter_core_core_fsm
module filter_core_core_fsm (
  clk, rst, fsm_output, buffer_buf_vinit_C_1_tr0
);
  input clk;
  input rst;
  output [6:0] fsm_output;
  reg [6:0] fsm_output;
  input buffer_buf_vinit_C_1_tr0;


  // FSM State Type Declaration for filter_core_core_fsm_1
  parameter
    core_rlp_C_0 = 3'd0,
    buffer_buf_vinit_C_0 = 3'd1,
    buffer_buf_vinit_C_1 = 3'd2,
    main_C_0 = 3'd3,
    main_C_1 = 3'd4,
    main_C_2 = 3'd5,
    main_C_3 = 3'd6;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : filter_core_core_fsm_1
    case (state_var)
      buffer_buf_vinit_C_0 : begin
        fsm_output = 7'b10;
        state_var_NS = buffer_buf_vinit_C_1;
      end
      buffer_buf_vinit_C_1 : begin
        fsm_output = 7'b100;
        if ( buffer_buf_vinit_C_1_tr0 ) begin
          state_var_NS = buffer_buf_vinit_C_0;
        end
        else begin
          state_var_NS = main_C_0;
        end
      end
      main_C_0 : begin
        fsm_output = 7'b1000;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 7'b10000;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 7'b100000;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 7'b1000000;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 7'b1;
        state_var_NS = buffer_buf_vinit_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule
`endif

// ------------------------------------------------------------------
//  Design Unit:    filter_core
// ------------------------------------------------------------------


`ifdef filter_core
`else
`define filter_core
module filter_core (
  clk, rst, in_data_rsc_z, in_data_rsc_lz, in_data_vld_rsc_z, out_data_rsc_z, out_data_rsc_lz,
      mcu_data_rsci_adr_d, mcu_data_rsci_d_d, mcu_data_rsci_we_d, mcu_data_rsci_q_d,
      mcu_data_rsci_ram_rw_A_internal_RMASK_B_d, buffer_buf_rsci_radr_d, buffer_buf_rsci_wadr_d,
      buffer_buf_rsci_d_d, buffer_buf_rsci_we_d, buffer_buf_rsci_re_d, buffer_buf_rsci_q_d
);
  input clk;
  input rst;
  input [2:0] in_data_rsc_z;
  output in_data_rsc_lz;
  input in_data_vld_rsc_z;
  output [2:0] out_data_rsc_z;
  output out_data_rsc_lz;
  output [8:0] mcu_data_rsci_adr_d;
  output [31:0] mcu_data_rsci_d_d;
  output mcu_data_rsci_we_d;
  input [31:0] mcu_data_rsci_q_d;
  output mcu_data_rsci_ram_rw_A_internal_RMASK_B_d;
  output [9:0] buffer_buf_rsci_radr_d;
  output [9:0] buffer_buf_rsci_wadr_d;
  output [2:0] buffer_buf_rsci_d_d;
  output buffer_buf_rsci_we_d;
  output buffer_buf_rsci_re_d;
  input [2:0] buffer_buf_rsci_q_d;


  // Interconnect Declarations
  reg in_data_rsci_ld;
  wire [2:0] in_data_rsci_d;
  wire in_data_vld_rsci_d;
  reg out_data_rsci_ld;
  reg out_data_rsci_d_0;
  wire [6:0] fsm_output;
  wire if_if_if_and_tmp;
  wire [2:0] pixel_processing_if_if_acc_tmp;
  wire [3:0] nl_pixel_processing_if_if_acc_tmp;
  wire clip_window_clip_window_nor_tmp;
  wire clip_window_clip_window_nor_1_tmp;
  wire system_input_system_input_or_tmp;
  wire clip_window_clip_window_and_1_tmp;
  wire clip_window_clip_window_and_tmp;
  wire and_2_tmp;
  wire system_input_system_input_nand_tmp;
  wire or_dcpl;
  wire and_dcpl_11;
  wire and_dcpl_33;
  wire and_dcpl_44;
  wire and_dcpl_45;
  wire and_dcpl_57;
  wire nor_tmp_4;
  wire mux_tmp_3;
  wire and_dcpl_64;
  wire or_tmp_33;
  wire or_tmp_42;
  wire or_tmp_48;
  wire or_tmp_56;
  reg mcu_ready_sva;
  reg [2:0] pixel_processing_threshold_sva;
  reg [8:0] pixel_processing_frame_sva;
  wire [9:0] nl_pixel_processing_frame_sva;
  reg [31:0] system_input_c_sva;
  reg [31:0] system_input_r_sva;
  reg [31:0] system_input_c_filter_sva;
  reg [31:0] system_input_r_filter_sva;
  reg system_input_output_vld_sva;
  reg [2:0] system_input_window_4_sva;
  reg [2:0] system_input_window_3_sva;
  reg [2:0] system_input_window_5_sva;
  reg [2:0] system_input_window_6_sva;
  reg [2:0] system_input_window_7_sva;
  reg [2:0] system_input_window_8_sva;
  reg [9:0] buffer_buf_vinit_ndx_sva;
  reg buffer_sel_1_0_sva_1;
  reg if_if_if_and_mdf_sva_2;
  reg else_io_read_in_data_vld_rsc_svs;
  reg [2:0] system_input_din_sva_1;
  reg buffer_sel_1_0_sva_dfm;
  reg [2:0] buffer_t0_sva_1;
  reg clip_window_first_row_0_sva_5;
  reg clip_window_last_row_0_sva_7;
  reg clip_window_last_col_0_sva_3;
  reg system_input_output_vld_sva_dfm;
  reg system_input_land_1_lpi_1_dfm_1;
  reg [2:0] median_max2_5_1_lpi_1_dfm;
  reg [2:0] median_max_4_2_lpi_1_dfm;
  reg [2:0] median_max2_3_2_lpi_1_dfm;
  reg [2:0] median_max_2_2_lpi_1_dfm;
  reg [2:0] median_max2_1_lpi_1_dfm;
  reg [2:0] median_max_4_1_lpi_1_dfm;
  reg [2:0] median_max_6_lpi_1_dfm;
  reg [2:0] median_max_5_3_lpi_1_dfm;
  reg [2:0] median_max_7_lpi_1_dfm;
  reg pixel_processing_if_if_1_pixel_processing_if_if_1_if_and_svs_1;
  reg buffer_buf_buffer_buf_nor_itm_1;
  reg [9:0] buffer_buf_acc_itm_2;
  wire [10:0] nl_buffer_buf_acc_itm_2;
  reg [2:0] median_max_5_lpi_1_dfm_5;
  reg asn_itm;
  reg else_io_read_in_data_vld_rsc_svs_st_1;
  reg [3:0] buffer_acc_1_itm_2;
  wire [4:0] nl_buffer_acc_1_itm_2;
  reg [3:0] buffer_acc_3_itm_2;
  wire [4:0] nl_buffer_acc_3_itm_2;
  reg [5:0] buffer_slc_buffer_c_5_0_1_itm_2;
  reg system_input_output_vld_sva_dfm_st_1;
  reg [2:0] clip_window_switch_lp_3_asn_2_itm;
  reg pixel_processing_if_pixel_processing_if_if_nor_itm;
  reg [2:0] pixel_processing_if_asn_itm;
  reg [8:0] pixel_processing_if_if_1_asn_itm;
  reg and_itm;
  reg asn_itm_1;
  reg else_io_read_in_data_vld_rsc_svs_st_2;
  reg system_input_output_vld_sva_dfm_st_2;
  reg pixel_processing_if_pixel_processing_if_if_nor_itm_2;
  reg main_stage_0_2;
  reg and_2_cse;
  wire and_116_cse;
  wire and_120_cse;
  wire and_128_cse;
  wire and_143_cse;
  wire and_146_cse;
  wire and_147_cse;
  wire and_148_cse;
  wire and_154_cse;
  wire and_141_cse;
  wire pixel_processing_if_if_1_pixel_processing_if_if_1_if_and_svs;
  wire system_input_land_1_lpi_1_dfm;
  wire [2:0] median_max_8_lpi_1_dfm_mx0;
  wire [2:0] median_max2_9_lpi_1_dfm_1_mx0;
  wire [2:0] median_max2_2_lpi_1_dfm_mx0;
  wire [2:0] pixel_processing_window_8_lpi_1_dfm;
  wire [2:0] pixel_processing_window_6_lpi_1_dfm;
  wire [2:0] median_max2_0_lpi_1_dfm_1_mx0;
  wire [2:0] median_max_1_2_lpi_1_dfm_mx0;
  wire [2:0] pixel_processing_window_2_lpi_1_dfm;
  wire [2:0] pixel_processing_window_0_lpi_1_dfm;
  wire [2:0] median_max_4_lpi_1_dfm_mx0;
  wire [2:0] median_max2_8_2_lpi_1_dfm_mx0;
  wire [2:0] median_max_3_lpi_1_dfm_mx0;
  wire [2:0] median_max2_5_2_lpi_1_dfm_mx0;
  wire [2:0] median_max2_9_lpi_1_dfm_mx0;
  wire [2:0] median_max2_4_2_lpi_1_dfm_mx0;
  wire [2:0] median_max_6_2_lpi_1_dfm_mx0;
  wire [2:0] median_max2_7_1_lpi_1_dfm_mx0;
  wire [2:0] median_max_5_2_lpi_1_dfm_mx0;
  wire [2:0] median_max2_6_1_lpi_1_dfm_mx0;
  wire [2:0] buffer_qr_1_lpi_1_dfm_mx0;
  wire [2:0] median_max2_0_lpi_1_dfm_mx0;
  wire [2:0] median_max_3_1_lpi_1_dfm_mx0;
  wire [2:0] median_max2_1_1_lpi_1_dfm_mx0;
  wire [2:0] median_max2_4_1_lpi_1_dfm_mx0;
  wire [2:0] clip_window_qr_lpi_1_dfm_mx0;
  wire [2:0] median_max2_6_2_lpi_1_dfm_mx0;
  wire [2:0] median_max2_7_2_lpi_1_dfm_mx0;
  wire [2:0] median_max_7_1_lpi_1_dfm_mx0;
  wire [2:0] median_max_8_1_lpi_1_dfm_mx0;
  wire [2:0] median_max2_8_1_lpi_1_dfm_mx0;
  wire [2:0] clip_window_qr_2_lpi_1_dfm_mx0;
  wire [2:0] median_max_1_1_lpi_1_dfm_mx0;
  wire [2:0] median_max_2_1_lpi_1_dfm_mx0;
  wire [2:0] median_max2_2_1_lpi_1_dfm_mx0;
  wire [2:0] median_max2_3_1_lpi_1_dfm_mx0;
  wire [2:0] clip_window_qr_3_lpi_1_dfm_mx0;
  wire reg_system_input_system_input_output_vld_and_cse;
  wire nand_2_cse;
  wire mcu_data_rsci_adr_d_mx0c2;
  wire mcu_data_rsci_adr_d_mx0c3;
  wire [2:0] median_max_5_lpi_1_dfm_mx0;
  wire L1a_if_slc_L1a_if_acc_14_3_itm;
  wire L1a_if_slc_L1a_if_acc_13_3_itm;
  wire L1a_if_slc_L1a_if_acc_12_3_itm;
  wire L1b_if_slc_L1b_if_acc_12_3_itm;
  wire L1b_if_slc_L1b_if_acc_11_3_itm;
  wire L1a_if_slc_L1a_if_acc_4_3_itm;
  wire [2:0] L1b_asn_4_mx1w1;
  wire [2:0] L1b_asn_44_mx0w1;
  wire buffer_sel_1_0_sva_dfm_mx0;
  wire [2:0] pixel_processing_if_if_acc_2_psp_sva;
  wire [3:0] nl_pixel_processing_if_if_acc_2_psp_sva;
  wire [2:0] pixel_processing_if_if_acc_8_psp;
  wire [3:0] nl_pixel_processing_if_if_acc_8_psp;
  wire [3:0] pixel_processing_if_if_acc_6_sdt;
  wire [4:0] nl_pixel_processing_if_if_acc_6_sdt;
  wire [2:0] median_max2_2_2_lpi_1_dfm_mx0;
  wire clip_window_switch_lp_equal_tmp;
  wire clip_window_switch_lp_equal_tmp_1;
  wire clip_window_switch_lp_equal_tmp_2;
  wire clip_window_switch_lp_2_equal_tmp;
  wire clip_window_switch_lp_2_equal_tmp_1;
  wire clip_window_switch_lp_2_equal_tmp_2;
  wire [2:0] median_max2_8_lpi_1_dfm_mx0;
  wire [2:0] L1a_asn_11_mx0w1;
  wire [2:0] median_max2_7_lpi_1_dfm_mx0;
  wire [2:0] L1a_asn_16_mx0w1;
  wire [2:0] median_max2_5_3_lpi_1_dfm_mx0;
  wire [2:0] median_max_2_lpi_1_dfm_mx0;
  wire [2:0] median_max2_4_lpi_1_dfm_mx0;
  wire [2:0] median_max_7_2_lpi_1_dfm_mx0;
  wire [2:0] median_max_5_1_lpi_1_dfm_mx0;
  wire clip_window_switch_lp_1_equal_tmp;
  wire clip_window_switch_lp_1_equal_tmp_1;
  wire clip_window_switch_lp_1_equal_tmp_2;
  wire [2:0] buffer_qr_lpi_1_dfm_mx0;
  wire clip_window_switch_lp_3_equal_tmp;
  wire clip_window_switch_lp_3_equal_tmp_1;
  wire clip_window_switch_lp_3_equal_tmp_2;
  wire [2:0] median_max2_6_lpi_1_dfm_mx0;
  wire [2:0] median_max2_5_lpi_1_dfm_mx0;
  wire L1b_if_acc_15_itm_3;
  wire L1b_if_acc_14_itm_3;
  wire L1b_if_acc_13_itm_3;
  wire and_104_rgt;
  wire median_max_and_7_rgt;
  wire and_108_rgt;
  wire reg_median_median_max_or_2_cse;
  wire reg_pixel_processing_if_pixel_processing_if_if_pixel_processing_if_if_and_cse;
  wire z_out_3;
  wire z_out_1_3;
  wire z_out_2_3;
  wire z_out_3_3;
  wire z_out_4_3;
  wire z_out_5_3;
  wire z_out_6_3;
  wire z_out_7_3;
  wire z_out_8_3;

  wire[31:0] system_input_if_2_qelse_acc_nl;
  wire[32:0] nl_system_input_if_2_qelse_acc_nl;
  wire[0:0] system_input_if_2_system_input_if_2_nand_nl;
  wire[31:0] system_input_if_1_qelse_acc_nl;
  wire[32:0] nl_system_input_if_1_qelse_acc_nl;
  wire[0:0] clip_window_switch_lp_2_not_4_nl;
  wire[31:0] system_input_else_2_acc_nl;
  wire[32:0] nl_system_input_else_2_acc_nl;
  wire[0:0] and_102_nl;
  wire[0:0] median_max2_and_5_nl;
  wire[0:0] median_max_and_3_nl;
  wire[0:0] median_max2_and_3_nl;
  wire[0:0] median_max_and_1_nl;
  wire[0:0] median_max2_median_max2_nor_nl;
  wire[0:0] buffer_nor_nl;
  wire[1:0] pixel_processing_if_if_acc_7_nl;
  wire[2:0] nl_pixel_processing_if_if_acc_7_nl;
  wire[2:0] pixel_processing_if_if_acc_5_nl;
  wire[3:0] nl_pixel_processing_if_if_acc_5_nl;
  wire[2:0] pixel_processing_if_if_acc_4_nl;
  wire[3:0] nl_pixel_processing_if_if_acc_4_nl;
  wire[0:0] nor_nl;
  wire[0:0] clip_window_switch_lp_2_nor_nl;
  wire[0:0] clip_window_switch_lp_nor_nl;
  wire[0:0] clip_window_switch_lp_3_nor_nl;
  wire[0:0] clip_window_switch_lp_1_nor_nl;
  wire[3:0] L1b_if_acc_15_nl;
  wire[5:0] nl_L1b_if_acc_15_nl;
  wire[3:0] L1b_if_acc_14_nl;
  wire[5:0] nl_L1b_if_acc_14_nl;
  wire[3:0] L1b_if_acc_13_nl;
  wire[5:0] nl_L1b_if_acc_13_nl;
  wire[0:0] nand_6_nl;
  wire[3:0] L1a_if_acc_14_nl;
  wire[5:0] nl_L1a_if_acc_14_nl;
  wire[3:0] L1a_if_acc_13_nl;
  wire[5:0] nl_L1a_if_acc_13_nl;
  wire[3:0] L1a_if_acc_12_nl;
  wire[5:0] nl_L1a_if_acc_12_nl;
  wire[3:0] L1b_if_acc_12_nl;
  wire[5:0] nl_L1b_if_acc_12_nl;
  wire[3:0] L1b_if_acc_11_nl;
  wire[5:0] nl_L1b_if_acc_11_nl;
  wire[3:0] L1a_if_acc_4_nl;
  wire[5:0] nl_L1a_if_acc_4_nl;
  wire[0:0] mcu_data_mcu_data_or_nl;
  wire[2:0] mcu_data_and_1_nl;
  wire[2:0] mcu_data_mux1h_1_nl;
  wire[0:0] mcu_data_nor_1_nl;
  wire[0:0] mux_56_nl;
  wire[0:0] mux_55_nl;
  wire[0:0] nand_1_nl;
  wire[31:0] mcu_data_mux1h_nl;
  wire[31:0] pixel_processing_if_if_pixel_processing_if_if_acc_1_nl;
  wire[32:0] nl_pixel_processing_if_if_pixel_processing_if_if_acc_1_nl;
  wire[0:0] mcu_data_nor_2_nl;
  wire[9:0] buffer_buf_mux_3_nl;
  wire[0:0] buffer_buf_nor_nl;
  wire[9:0] buffer_buf_mux_2_nl;
  wire[0:0] buffer_buf_nor_1_nl;
  wire[4:0] acc_nl;
  wire[5:0] nl_acc_nl;
  wire[2:0] thresholding_if_mux1h_3_nl;
  wire[2:0] thresholding_if_mux1h_4_nl;
  wire[4:0] acc_1_nl;
  wire[5:0] nl_acc_1_nl;
  wire[2:0] L1b_if_mux1h_3_nl;
  wire[2:0] L1b_if_mux1h_4_nl;
  wire[4:0] acc_2_nl;
  wire[5:0] nl_acc_2_nl;
  wire[2:0] L1a_if_mux1h_6_nl;
  wire[2:0] L1a_if_mux1h_7_nl;
  wire[2:0] clip_window_mux_2_nl;
  wire[4:0] acc_3_nl;
  wire[5:0] nl_acc_3_nl;
  wire[2:0] L1a_if_mux1h_8_nl;
  wire[2:0] L1a_if_mux1h_9_nl;
  wire[4:0] acc_4_nl;
  wire[5:0] nl_acc_4_nl;
  wire[2:0] L1a_if_mux_9_nl;
  wire[2:0] L1a_if_mux_10_nl;
  wire[4:0] acc_5_nl;
  wire[5:0] nl_acc_5_nl;
  wire[2:0] L1a_if_mux_11_nl;
  wire[2:0] L1a_if_mux_12_nl;
  wire[4:0] acc_6_nl;
  wire[5:0] nl_acc_6_nl;
  wire[2:0] L1b_if_mux_6_nl;
  wire[2:0] L1b_if_mux_7_nl;
  wire[4:0] acc_7_nl;
  wire[5:0] nl_acc_7_nl;
  wire[2:0] L1a_if_mux_13_nl;
  wire[2:0] L1a_if_mux_14_nl;
  wire[4:0] acc_8_nl;
  wire[5:0] nl_acc_8_nl;
  wire[2:0] L1b_if_mux_8_nl;
  wire[2:0] L1b_if_mux_9_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [2:0] nl_out_data_rsci_d;
  assign nl_out_data_rsci_d = {{2{out_data_rsci_d_0}}, out_data_rsci_d_0};
  wire [0:0] nl_filter_core_core_fsm_inst_buffer_buf_vinit_C_1_tr0;
  assign nl_filter_core_core_fsm_inst_buffer_buf_vinit_C_1_tr0 = ~ buffer_buf_buffer_buf_nor_itm_1;
  mgc_in_wire_en_v1 #(.rscid(32'sd1),
  .width(32'sd3)) in_data_rsci (
      .ld(in_data_rsci_ld),
      .d(in_data_rsci_d),
      .lz(in_data_rsc_lz),
      .z(in_data_rsc_z)
    );
  mgc_in_wire_v1 #(.rscid(32'sd2),
  .width(32'sd1)) in_data_vld_rsci (
      .d(in_data_vld_rsci_d),
      .z(in_data_vld_rsc_z)
    );
  mgc_out_stdreg_en_v1 #(.rscid(32'sd3),
  .width(32'sd3)) out_data_rsci (
      .ld(out_data_rsci_ld),
      .d(nl_out_data_rsci_d[2:0]),
      .lz(out_data_rsc_lz),
      .z(out_data_rsc_z)
    );
  filter_core_core_fsm filter_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .buffer_buf_vinit_C_1_tr0(nl_filter_core_core_fsm_inst_buffer_buf_vinit_C_1_tr0[0:0])
    );
  assign reg_system_input_system_input_output_vld_and_cse = in_data_vld_rsci_d &
      mcu_ready_sva & (fsm_output[3]);
  assign reg_pixel_processing_if_pixel_processing_if_if_pixel_processing_if_if_and_cse
      = mcu_ready_sva & (~ or_tmp_56);
  assign and_104_rgt = mcu_ready_sva & (~ L1b_if_acc_15_itm_3) & (fsm_output[5]);
  assign median_max_and_7_rgt = mcu_ready_sva & (~ L1b_if_acc_14_itm_3) & (fsm_output[5]);
  assign reg_median_median_max_or_2_cse = (mcu_ready_sva & L1b_if_acc_14_itm_3 &
      (fsm_output[5])) | median_max_and_7_rgt;
  assign and_108_rgt = mcu_ready_sva & (~ L1b_if_acc_13_itm_3) & (fsm_output[5]);
  assign L1b_asn_4_mx1w1 = MUX_v_3_2_2(median_max_7_2_lpi_1_dfm_mx0, L1a_asn_11_mx0w1,
      L1a_if_slc_L1a_if_acc_14_3_itm);
  assign median_max_5_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_6_lpi_1_dfm_mx0, median_max2_5_lpi_1_dfm_mx0,
      z_out_1_3);
  assign system_input_system_input_or_tmp = system_input_output_vld_sva | ((system_input_c_sva==32'b00000000000000000000000000000001)
      & (system_input_r_sva==32'b00000000000000000000000000000001));
  assign clip_window_clip_window_and_tmp = (system_input_r_filter_sva==32'b00000000000000000000000011101111);
  assign pixel_processing_if_if_1_pixel_processing_if_if_1_if_and_svs = (pixel_processing_frame_sva[0])
      & (pixel_processing_if_if_acc_tmp==3'b000);
  assign system_input_land_1_lpi_1_dfm = clip_window_clip_window_and_1_tmp & clip_window_clip_window_and_tmp;
  assign L1b_asn_44_mx0w1 = MUX_v_3_2_2(median_max2_0_lpi_1_dfm_mx0, median_max_1_1_lpi_1_dfm_mx0,
      z_out_7_3);
  assign clip_window_clip_window_nor_tmp = ~((system_input_r_filter_sva!=32'b00000000000000000000000000000000));
  assign clip_window_clip_window_and_1_tmp = (system_input_c_filter_sva==32'b00000000000000000000000100111111);
  assign buffer_nor_nl = ~((system_input_c_sva!=32'b00000000000000000000000000000000));
  assign buffer_sel_1_0_sva_dfm_mx0 = MUX_s_1_2_2(buffer_sel_1_0_sva_1, (~ buffer_sel_1_0_sva_1),
      buffer_nor_nl);
  assign nl_pixel_processing_if_if_acc_tmp = conv_u2u_1_3(pixel_processing_if_if_acc_2_psp_sva[2])
      + conv_u2u_2_3(pixel_processing_if_if_acc_2_psp_sva[1:0]);
  assign pixel_processing_if_if_acc_tmp = nl_pixel_processing_if_if_acc_tmp[2:0];
  assign nl_pixel_processing_if_if_acc_7_nl = conv_s2s_1_2(~ (pixel_processing_if_if_acc_8_psp[2]))
      + conv_u2s_1_2(~ (pixel_processing_if_if_acc_8_psp[1]));
  assign pixel_processing_if_if_acc_7_nl = nl_pixel_processing_if_if_acc_7_nl[1:0];
  assign nl_pixel_processing_if_if_acc_2_psp_sva = conv_s2u_2_3(pixel_processing_if_if_acc_7_nl)
      + ({(pixel_processing_if_if_acc_8_psp[2]) , (pixel_processing_if_if_acc_8_psp[0])
      , (pixel_processing_if_if_acc_6_sdt[0])});
  assign pixel_processing_if_if_acc_2_psp_sva = nl_pixel_processing_if_if_acc_2_psp_sva[2:0];
  assign nl_pixel_processing_if_if_acc_8_psp = (pixel_processing_if_if_acc_6_sdt[3:1])
      + 3'b101;
  assign pixel_processing_if_if_acc_8_psp = nl_pixel_processing_if_if_acc_8_psp[2:0];
  assign nl_pixel_processing_if_if_acc_5_nl = conv_u2u_2_3(pixel_processing_frame_sva[2:1])
      + conv_u2u_2_3(~ (pixel_processing_frame_sva[4:3]));
  assign pixel_processing_if_if_acc_5_nl = nl_pixel_processing_if_if_acc_5_nl[2:0];
  assign nl_pixel_processing_if_if_acc_4_nl = conv_u2u_2_3(pixel_processing_frame_sva[6:5])
      + conv_u2u_2_3(~ (pixel_processing_frame_sva[8:7]));
  assign pixel_processing_if_if_acc_4_nl = nl_pixel_processing_if_if_acc_4_nl[2:0];
  assign nl_pixel_processing_if_if_acc_6_sdt = conv_u2u_3_4(pixel_processing_if_if_acc_5_nl)
      + conv_u2u_3_4(pixel_processing_if_if_acc_4_nl);
  assign pixel_processing_if_if_acc_6_sdt = nl_pixel_processing_if_if_acc_6_sdt[3:0];
  assign median_max2_0_lpi_1_dfm_1_mx0 = MUX_v_3_2_2(median_max_1_1_lpi_1_dfm_mx0,
      median_max2_0_lpi_1_dfm_mx0, z_out_7_3);
  assign median_max_1_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_2_2_lpi_1_dfm_mx0,
      L1b_asn_44_mx0w1, z_out_1_3);
  assign median_max2_2_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_3_1_lpi_1_dfm_mx0,
      median_max_2_1_lpi_1_dfm_mx0, z_out_5_3);
  assign median_max_2_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_1_1_lpi_1_dfm_mx0,
      median_max2_2_1_lpi_1_dfm_mx0, z_out_8_3);
  assign median_max_3_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_4_1_lpi_1_dfm_mx0,
      median_max2_3_1_lpi_1_dfm_mx0, z_out_6_3);
  assign median_max2_0_lpi_1_dfm_mx0 = MUX_v_3_2_2(clip_window_qr_lpi_1_dfm_mx0,
      pixel_processing_window_0_lpi_1_dfm, z_out_3_3);
  assign median_max_1_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_2_1_lpi_1_dfm_mx0,
      median_max2_1_1_lpi_1_dfm_mx0, z_out_8_3);
  assign median_max2_3_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(pixel_processing_window_2_lpi_1_dfm,
      clip_window_qr_3_lpi_1_dfm_mx0, z_out_4_3);
  assign nor_nl = ~(clip_window_clip_window_and_tmp | z_out_2_3);
  assign median_max2_4_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(system_input_window_7_sva, system_input_window_8_sva,
      nor_nl);
  assign median_max2_1_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(pixel_processing_window_0_lpi_1_dfm,
      clip_window_qr_lpi_1_dfm_mx0, z_out_3_3);
  assign median_max2_2_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(clip_window_qr_3_lpi_1_dfm_mx0,
      pixel_processing_window_2_lpi_1_dfm, z_out_4_3);
  assign clip_window_switch_lp_2_nor_nl = ~(clip_window_switch_lp_2_equal_tmp | clip_window_switch_lp_2_equal_tmp_1
      | clip_window_switch_lp_2_equal_tmp_2);
  assign pixel_processing_window_2_lpi_1_dfm = MUX1HOT_v_3_4_2(system_input_window_7_sva,
      system_input_window_4_sva, system_input_window_8_sva, system_input_window_5_sva,
      {(clip_window_switch_lp_2_nor_nl) , clip_window_switch_lp_2_equal_tmp , clip_window_switch_lp_2_equal_tmp_1
      , clip_window_switch_lp_2_equal_tmp_2});
  assign clip_window_qr_3_lpi_1_dfm_mx0 = MUX_v_3_2_2(system_input_window_6_sva,
      system_input_window_7_sva, clip_window_clip_window_nor_tmp);
  assign clip_window_switch_lp_nor_nl = ~(clip_window_switch_lp_equal_tmp | clip_window_switch_lp_equal_tmp_1
      | clip_window_switch_lp_equal_tmp_2);
  assign pixel_processing_window_0_lpi_1_dfm = MUX1HOT_v_3_4_2(system_input_window_7_sva,
      system_input_window_4_sva, system_input_window_6_sva, system_input_window_3_sva,
      {(clip_window_switch_lp_nor_nl) , clip_window_switch_lp_equal_tmp , clip_window_switch_lp_equal_tmp_1
      , clip_window_switch_lp_equal_tmp_2});
  assign clip_window_qr_lpi_1_dfm_mx0 = MUX_v_3_2_2(system_input_window_4_sva, system_input_window_7_sva,
      clip_window_clip_window_nor_1_tmp);
  assign clip_window_clip_window_nor_1_tmp = ~((system_input_c_filter_sva!=32'b00000000000000000000000000000000));
  assign clip_window_switch_lp_equal_tmp = clip_window_clip_window_nor_tmp & (~ clip_window_clip_window_nor_1_tmp);
  assign clip_window_switch_lp_equal_tmp_1 = clip_window_clip_window_nor_1_tmp &
      (~ clip_window_clip_window_nor_tmp);
  assign clip_window_switch_lp_equal_tmp_2 = ~(clip_window_clip_window_nor_1_tmp
      | clip_window_clip_window_nor_tmp);
  assign clip_window_switch_lp_2_equal_tmp = clip_window_clip_window_and_tmp & (~
      clip_window_clip_window_nor_1_tmp);
  assign clip_window_switch_lp_2_equal_tmp_1 = clip_window_clip_window_nor_1_tmp
      & (~ clip_window_clip_window_and_tmp);
  assign clip_window_switch_lp_2_equal_tmp_2 = ~(clip_window_clip_window_nor_1_tmp
      | clip_window_clip_window_and_tmp);
  assign system_input_system_input_nand_tmp = ~((system_input_c_sva==32'b00000000000000000000000100111111));
  assign and_2_tmp = in_data_vld_rsci_d & mcu_ready_sva;
  assign if_if_if_and_tmp = (mcu_data_rsci_q_d==32'b00000000000000000000000000000001);
  assign median_max2_8_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_9_lpi_1_dfm_1_mx0,
      median_max_8_lpi_1_dfm_mx0, z_out_3);
  assign L1a_asn_11_mx0w1 = MUX_v_3_2_2(median_max_4_lpi_1_dfm_mx0, median_max2_6_2_lpi_1_dfm_mx0,
      L1b_if_slc_L1b_if_acc_11_3_itm);
  assign median_max2_7_lpi_1_dfm_mx0 = MUX_v_3_2_2(L1a_asn_11_mx0w1, median_max_7_2_lpi_1_dfm_mx0,
      L1a_if_slc_L1a_if_acc_14_3_itm);
  assign L1a_asn_16_mx0w1 = MUX_v_3_2_2(median_max_2_2_lpi_1_dfm, median_max_3_lpi_1_dfm_mx0,
      z_out_7_3);
  assign median_max2_5_3_lpi_1_dfm_mx0 = MUX_v_3_2_2(L1a_asn_16_mx0w1, median_max_5_1_lpi_1_dfm_mx0,
      L1a_if_slc_L1a_if_acc_13_3_itm);
  assign median_max_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_1_lpi_1_dfm, median_max2_2_lpi_1_dfm_mx0,
      z_out_1_3);
  assign median_max2_4_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_5_1_lpi_1_dfm_mx0,
      L1a_asn_16_mx0w1, L1a_if_slc_L1a_if_acc_13_3_itm);
  assign median_max2_9_lpi_1_dfm_1_mx0 = MUX_v_3_2_2(median_max_8_1_lpi_1_dfm_mx0,
      median_max2_9_lpi_1_dfm_mx0, L1a_if_slc_L1a_if_acc_12_3_itm);
  assign median_max_8_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_7_2_lpi_1_dfm_mx0,
      median_max2_8_2_lpi_1_dfm_mx0, L1b_if_slc_L1b_if_acc_12_3_itm);
  assign median_max_7_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_8_2_lpi_1_dfm_mx0,
      median_max2_7_2_lpi_1_dfm_mx0, L1b_if_slc_L1b_if_acc_12_3_itm);
  assign median_max_5_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_6_2_lpi_1_dfm_mx0,
      median_max_4_lpi_1_dfm_mx0, L1b_if_slc_L1b_if_acc_11_3_itm);
  assign median_max2_8_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_9_lpi_1_dfm_mx0,
      median_max_8_1_lpi_1_dfm_mx0, L1a_if_slc_L1a_if_acc_12_3_itm);
  assign median_max2_7_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_5_2_lpi_1_dfm_mx0,
      median_max_7_1_lpi_1_dfm_mx0, z_out_5_3);
  assign median_max_4_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_3_2_lpi_1_dfm, median_max2_4_2_lpi_1_dfm_mx0,
      z_out_6_3);
  assign median_max2_6_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_7_1_lpi_1_dfm_mx0,
      median_max2_5_2_lpi_1_dfm_mx0, z_out_5_3);
  assign median_max2_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_3_lpi_1_dfm_mx0, median_max_2_2_lpi_1_dfm,
      z_out_7_3);
  assign median_max2_9_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_7_1_lpi_1_dfm_mx0,
      pixel_processing_window_8_lpi_1_dfm, z_out_2_3);
  assign median_max_8_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_6_2_lpi_1_dfm_mx0,
      median_max2_8_1_lpi_1_dfm_mx0, z_out_8_3);
  assign median_max2_5_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_4_2_lpi_1_dfm, median_max_5_2_lpi_1_dfm_mx0,
      z_out_3_3);
  assign median_max_7_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_8_1_lpi_1_dfm_mx0,
      median_max_6_2_lpi_1_dfm_mx0, z_out_8_3);
  assign median_max_3_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_4_2_lpi_1_dfm_mx0,
      median_max2_3_2_lpi_1_dfm, z_out_6_3);
  assign median_max_6_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_5_1_lpi_1_dfm, median_max2_6_1_lpi_1_dfm_mx0,
      z_out_4_3);
  assign median_max2_8_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(pixel_processing_window_8_lpi_1_dfm,
      median_max2_7_1_lpi_1_dfm_mx0, z_out_2_3);
  assign median_max2_4_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_5_2_lpi_1_dfm_mx0,
      median_max_4_2_lpi_1_dfm, z_out_3_3);
  assign clip_window_switch_lp_3_nor_nl = ~(clip_window_switch_lp_3_equal_tmp | clip_window_switch_lp_3_equal_tmp_1
      | clip_window_switch_lp_3_equal_tmp_2);
  assign pixel_processing_window_8_lpi_1_dfm = MUX1HOT_v_3_4_2(system_input_window_7_sva,
      buffer_qr_1_lpi_1_dfm_mx0, clip_window_switch_lp_3_asn_2_itm, system_input_din_sva_1,
      {(clip_window_switch_lp_3_nor_nl) , clip_window_switch_lp_3_equal_tmp , clip_window_switch_lp_3_equal_tmp_1
      , clip_window_switch_lp_3_equal_tmp_2});
  assign median_max2_7_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(pixel_processing_window_6_lpi_1_dfm,
      clip_window_qr_2_lpi_1_dfm_mx0, L1a_if_slc_L1a_if_acc_4_3_itm);
  assign median_max_5_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_6_1_lpi_1_dfm_mx0,
      median_max2_5_1_lpi_1_dfm, z_out_4_3);
  assign median_max2_6_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(clip_window_qr_2_lpi_1_dfm_mx0,
      pixel_processing_window_6_lpi_1_dfm, L1a_if_slc_L1a_if_acc_4_3_itm);
  assign clip_window_switch_lp_1_nor_nl = ~(clip_window_switch_lp_1_equal_tmp | clip_window_switch_lp_1_equal_tmp_1
      | clip_window_switch_lp_1_equal_tmp_2);
  assign pixel_processing_window_6_lpi_1_dfm = MUX1HOT_v_3_4_2(system_input_window_7_sva,
      buffer_qr_1_lpi_1_dfm_mx0, system_input_window_6_sva, buffer_qr_lpi_1_dfm_mx0,
      {(clip_window_switch_lp_1_nor_nl) , clip_window_switch_lp_1_equal_tmp , clip_window_switch_lp_1_equal_tmp_1
      , clip_window_switch_lp_1_equal_tmp_2});
  assign clip_window_qr_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(buffer_qr_1_lpi_1_dfm_mx0,
      system_input_window_7_sva, clip_window_last_col_0_sva_3);
  assign buffer_qr_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(buffer_buf_rsci_q_d, buffer_t0_sva_1,
      buffer_sel_1_0_sva_dfm);
  assign clip_window_switch_lp_1_equal_tmp = clip_window_first_row_0_sva_5 & (~ clip_window_last_col_0_sva_3);
  assign clip_window_switch_lp_1_equal_tmp_1 = clip_window_last_col_0_sva_3 & (~
      clip_window_first_row_0_sva_5);
  assign clip_window_switch_lp_1_equal_tmp_2 = ~(clip_window_last_col_0_sva_3 | clip_window_first_row_0_sva_5);
  assign buffer_qr_lpi_1_dfm_mx0 = MUX_v_3_2_2(buffer_t0_sva_1, buffer_buf_rsci_q_d,
      buffer_sel_1_0_sva_dfm);
  assign clip_window_switch_lp_3_equal_tmp = clip_window_last_row_0_sva_7 & (~ clip_window_last_col_0_sva_3);
  assign clip_window_switch_lp_3_equal_tmp_1 = clip_window_last_col_0_sva_3 & (~
      clip_window_last_row_0_sva_7);
  assign clip_window_switch_lp_3_equal_tmp_2 = ~(clip_window_last_col_0_sva_3 | clip_window_last_row_0_sva_7);
  assign median_max2_6_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_7_lpi_1_dfm, median_max_6_lpi_1_dfm,
      z_out_2_3);
  assign median_max2_5_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_4_1_lpi_1_dfm, median_max_5_3_lpi_1_dfm,
      z_out_3_3);
  assign nl_L1b_if_acc_15_nl = ({1'b1 , median_max2_7_lpi_1_dfm_mx0}) + conv_u2u_3_4(~
      median_max2_8_lpi_1_dfm_mx0) + 4'b1;
  assign L1b_if_acc_15_nl = nl_L1b_if_acc_15_nl[3:0];
  assign L1b_if_acc_15_itm_3 = readslicef_4_1_3((L1b_if_acc_15_nl));
  assign nl_L1b_if_acc_14_nl = ({1'b1 , median_max2_5_3_lpi_1_dfm_mx0}) + conv_u2u_3_4(~
      L1b_asn_4_mx1w1) + 4'b1;
  assign L1b_if_acc_14_nl = nl_L1b_if_acc_14_nl[3:0];
  assign L1b_if_acc_14_itm_3 = readslicef_4_1_3((L1b_if_acc_14_nl));
  assign nl_L1b_if_acc_13_nl = ({1'b1 , median_max_2_lpi_1_dfm_mx0}) + conv_u2u_3_4(~
      median_max2_4_lpi_1_dfm_mx0) + 4'b1;
  assign L1b_if_acc_13_nl = nl_L1b_if_acc_13_nl[3:0];
  assign L1b_if_acc_13_itm_3 = readslicef_4_1_3((L1b_if_acc_13_nl));
  assign or_dcpl = ~(mcu_ready_sva & in_data_vld_rsci_d);
  assign and_dcpl_11 = else_io_read_in_data_vld_rsc_svs & system_input_output_vld_sva_dfm;
  assign and_dcpl_33 = mcu_ready_sva & else_io_read_in_data_vld_rsc_svs;
  assign and_dcpl_44 = asn_itm & else_io_read_in_data_vld_rsc_svs;
  assign and_dcpl_45 = and_dcpl_44 & system_input_output_vld_sva_dfm;
  assign and_dcpl_57 = system_input_land_1_lpi_1_dfm_1 & pixel_processing_if_if_1_pixel_processing_if_if_1_if_and_svs_1;
  assign nor_tmp_4 = system_input_land_1_lpi_1_dfm_1 & system_input_output_vld_sva_dfm
      & else_io_read_in_data_vld_rsc_svs & mcu_ready_sva;
  assign nand_6_nl = ~((~(system_input_land_1_lpi_1_dfm_1 & system_input_output_vld_sva_dfm
      & else_io_read_in_data_vld_rsc_svs)) & mcu_ready_sva);
  assign mux_tmp_3 = MUX_s_1_2_2(nor_tmp_4, (nand_6_nl), if_if_if_and_tmp);
  assign and_dcpl_64 = (~ asn_itm) & if_if_if_and_mdf_sva_2;
  assign nl_L1a_if_acc_14_nl = ({1'b1 , L1a_asn_11_mx0w1}) + conv_u2u_3_4(~ median_max_7_2_lpi_1_dfm_mx0)
      + 4'b1;
  assign L1a_if_acc_14_nl = nl_L1a_if_acc_14_nl[3:0];
  assign L1a_if_slc_L1a_if_acc_14_3_itm = readslicef_4_1_3((L1a_if_acc_14_nl));
  assign nl_L1a_if_acc_13_nl = ({1'b1 , L1a_asn_16_mx0w1}) + conv_u2u_3_4(~ median_max_5_1_lpi_1_dfm_mx0)
      + 4'b1;
  assign L1a_if_acc_13_nl = nl_L1a_if_acc_13_nl[3:0];
  assign L1a_if_slc_L1a_if_acc_13_3_itm = readslicef_4_1_3((L1a_if_acc_13_nl));
  assign nl_L1a_if_acc_12_nl = ({1'b1 , median_max_8_1_lpi_1_dfm_mx0}) + conv_u2u_3_4(~
      median_max2_9_lpi_1_dfm_mx0) + 4'b1;
  assign L1a_if_acc_12_nl = nl_L1a_if_acc_12_nl[3:0];
  assign L1a_if_slc_L1a_if_acc_12_3_itm = readslicef_4_1_3((L1a_if_acc_12_nl));
  assign nl_L1b_if_acc_12_nl = ({1'b1 , median_max2_7_2_lpi_1_dfm_mx0}) + conv_u2u_3_4(~
      median_max2_8_2_lpi_1_dfm_mx0) + 4'b1;
  assign L1b_if_acc_12_nl = nl_L1b_if_acc_12_nl[3:0];
  assign L1b_if_slc_L1b_if_acc_12_3_itm = readslicef_4_1_3((L1b_if_acc_12_nl));
  assign nl_L1b_if_acc_11_nl = ({1'b1 , median_max_4_lpi_1_dfm_mx0}) + conv_u2u_3_4(~
      median_max2_6_2_lpi_1_dfm_mx0) + 4'b1;
  assign L1b_if_acc_11_nl = nl_L1b_if_acc_11_nl[3:0];
  assign L1b_if_slc_L1b_if_acc_11_3_itm = readslicef_4_1_3((L1b_if_acc_11_nl));
  assign nl_L1a_if_acc_4_nl = ({1'b1 , pixel_processing_window_6_lpi_1_dfm}) + conv_u2u_3_4(~
      clip_window_qr_2_lpi_1_dfm_mx0) + 4'b1;
  assign L1a_if_acc_4_nl = nl_L1a_if_acc_4_nl[3:0];
  assign L1a_if_slc_L1a_if_acc_4_3_itm = readslicef_4_1_3((L1a_if_acc_4_nl));
  assign and_116_cse = and_2_tmp & (fsm_output[3]);
  assign and_120_cse = and_dcpl_33 & (fsm_output[4]);
  assign and_128_cse = (~(mcu_ready_sva & else_io_read_in_data_vld_rsc_svs)) & (fsm_output[4]);
  assign and_141_cse = and_dcpl_44 & system_input_output_vld_sva_dfm & pixel_processing_if_pixel_processing_if_if_nor_itm
      & (fsm_output[6]);
  assign and_143_cse = pixel_processing_if_pixel_processing_if_if_nor_itm_2 & system_input_output_vld_sva_dfm_st_2
      & else_io_read_in_data_vld_rsc_svs_st_2 & asn_itm_1 & main_stage_0_2 & (fsm_output[3]);
  assign and_146_cse = and_dcpl_64 & (fsm_output[6]);
  assign and_147_cse = ((~(pixel_processing_if_pixel_processing_if_if_nor_itm_2 &
      system_input_output_vld_sva_dfm_st_2 & else_io_read_in_data_vld_rsc_svs_st_2))
      | (~(asn_itm_1 & main_stage_0_2))) & (fsm_output[3]);
  assign and_148_cse = (~ mux_tmp_3) & (fsm_output[5]);
  assign and_154_cse = (~ mcu_ready_sva) & if_if_if_and_tmp & (fsm_output[5]);
  assign or_tmp_33 = nor_tmp_4 & (fsm_output[5]);
  assign or_tmp_42 = and_2_cse & (fsm_output[5]);
  assign or_tmp_48 = or_dcpl | (~ (fsm_output[3]));
  assign or_tmp_56 = (fsm_output[5:4]!=2'b00);
  assign mcu_data_rsci_adr_d_mx0c2 = and_154_cse | ((~ mcu_ready_sva) & (fsm_output[4]));
  assign mcu_data_rsci_adr_d_mx0c3 = and_146_cse | (and_dcpl_33 & system_input_output_vld_sva_dfm
      & and_dcpl_57 & (fsm_output[4]));
  assign nand_2_cse = ~(system_input_output_vld_sva_dfm & else_io_read_in_data_vld_rsc_svs);
  assign mcu_data_mcu_data_or_nl = mcu_data_rsci_adr_d_mx0c2 | mcu_data_rsci_adr_d_mx0c3
      | or_tmp_33;
  assign mcu_data_mux1h_1_nl = MUX1HOT_v_3_4_2(median_max_5_lpi_1_dfm_5, 3'b1, 3'b10,
      median_max_5_lpi_1_dfm_mx0, {and_143_cse , mcu_data_rsci_adr_d_mx0c3 , or_tmp_33
      , and_141_cse});
  assign nand_1_nl = ~(nand_2_cse & asn_itm);
  assign mux_55_nl = MUX_s_1_2_2(and_dcpl_45, (nand_1_nl), if_if_if_and_mdf_sva_2);
  assign mux_56_nl = MUX_s_1_2_2(and_dcpl_64, (mux_55_nl), pixel_processing_if_pixel_processing_if_if_nor_itm);
  assign mcu_data_nor_1_nl = ~(and_147_cse | and_148_cse | (fsm_output[2:0]!=3'b000)
      | ((~ (mux_56_nl)) & (fsm_output[6])) | ((nand_2_cse | (~(system_input_land_1_lpi_1_dfm_1
      & pixel_processing_if_if_1_pixel_processing_if_if_1_if_and_svs_1))) & mcu_ready_sva
      & (fsm_output[4])) | mcu_data_rsci_adr_d_mx0c2);
  assign mcu_data_and_1_nl = MUX_v_3_2_2(3'b000, (mcu_data_mux1h_1_nl), (mcu_data_nor_1_nl));
  assign mcu_data_rsci_adr_d = {5'b0 , (mcu_data_mcu_data_or_nl) , (mcu_data_and_1_nl)};
  assign nl_pixel_processing_if_if_pixel_processing_if_if_acc_1_nl = mcu_data_rsci_q_d
      + 32'b1;
  assign pixel_processing_if_if_pixel_processing_if_if_acc_1_nl = nl_pixel_processing_if_if_pixel_processing_if_if_acc_1_nl[31:0];
  assign mcu_data_mux1h_nl = MUX1HOT_v_32_4_2((pixel_processing_if_if_pixel_processing_if_if_acc_1_nl),
      32'b10, ({23'b0 , pixel_processing_if_if_1_asn_itm}), 32'b100, {and_143_cse
      , and_154_cse , or_tmp_33 , and_146_cse});
  assign mcu_data_nor_2_nl = ~(and_147_cse | and_148_cse | (~((fsm_output[6]) | (fsm_output[3])
      | (fsm_output[5]))) | ((asn_itm | (~ if_if_if_and_mdf_sva_2)) & (fsm_output[6])));
  assign mcu_data_rsci_d_d = MUX_v_32_2_2(32'b00000000000000000000000000000000, (mcu_data_mux1h_nl),
      (mcu_data_nor_2_nl));
  assign mcu_data_rsci_we_d = and_143_cse | (mux_tmp_3 & (fsm_output[5])) | and_146_cse;
  assign mcu_data_rsci_ram_rw_A_internal_RMASK_B_d = and_141_cse | ((~((~(and_dcpl_11
      & and_dcpl_57)) & mcu_ready_sva)) & (fsm_output[4]));
  assign buffer_buf_mux_3_nl = MUX_v_10_2_2((system_input_c_sva[9:0]), ({buffer_acc_1_itm_2
      , buffer_slc_buffer_c_5_0_1_itm_2}), and_120_cse);
  assign buffer_buf_nor_nl = ~((or_dcpl & (fsm_output[3])) | (~((fsm_output[4:3]!=2'b00)))
      | and_128_cse);
  assign buffer_buf_rsci_radr_d = MUX_v_10_2_2(10'b0000000000, (buffer_buf_mux_3_nl),
      (buffer_buf_nor_nl));
  assign buffer_buf_mux_2_nl = MUX_v_10_2_2(buffer_buf_vinit_ndx_sva, ({buffer_acc_3_itm_2
      , buffer_slc_buffer_c_5_0_1_itm_2}), and_120_cse);
  assign buffer_buf_nor_1_nl = ~((~((fsm_output[1]) | (fsm_output[4]))) | and_128_cse);
  assign buffer_buf_rsci_wadr_d = MUX_v_10_2_2(10'b0000000000, (buffer_buf_mux_2_nl),
      (buffer_buf_nor_1_nl));
  assign buffer_buf_rsci_d_d = MUX_v_3_2_2(3'b000, in_data_rsci_d, and_120_cse);
  assign buffer_buf_rsci_we_d = (fsm_output[1]) | and_120_cse;
  assign buffer_buf_rsci_re_d = and_116_cse | and_120_cse;
  always @(posedge clk) begin
    if ( rst ) begin
      out_data_rsci_d_0 <= 1'b0;
    end
    else if ( (fsm_output[6]) & asn_itm & else_io_read_in_data_vld_rsc_svs & system_input_output_vld_sva_dfm
        ) begin
      out_data_rsci_d_0 <= ~ z_out_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      out_data_rsci_ld <= 1'b0;
      in_data_rsci_ld <= 1'b0;
      buffer_buf_buffer_buf_nor_itm_1 <= 1'b0;
      buffer_buf_acc_itm_2 <= 10'b0;
      median_max_5_lpi_1_dfm_5 <= 3'b0;
      pixel_processing_if_pixel_processing_if_if_nor_itm_2 <= 1'b0;
      system_input_output_vld_sva_dfm_st_2 <= 1'b0;
      else_io_read_in_data_vld_rsc_svs_st_2 <= 1'b0;
      asn_itm_1 <= 1'b0;
      main_stage_0_2 <= 1'b0;
      buffer_slc_buffer_c_5_0_1_itm_2 <= 6'b0;
      buffer_acc_3_itm_2 <= 4'b0;
      buffer_acc_1_itm_2 <= 4'b0;
      else_io_read_in_data_vld_rsc_svs <= 1'b0;
      clip_window_switch_lp_3_asn_2_itm <= 3'b0;
      system_input_din_sva_1 <= 3'b0;
      buffer_t0_sva_1 <= 3'b0;
      if_if_if_and_mdf_sva_2 <= 1'b0;
    end
    else begin
      out_data_rsci_ld <= and_dcpl_45 & (fsm_output[6]);
      in_data_rsci_ld <= and_116_cse;
      buffer_buf_buffer_buf_nor_itm_1 <= ~((buffer_buf_vinit_ndx_sva!=10'b0000000000));
      buffer_buf_acc_itm_2 <= nl_buffer_buf_acc_itm_2[9:0];
      median_max_5_lpi_1_dfm_5 <= MUX_v_3_2_2(median_max2_5_lpi_1_dfm_mx0, median_max2_6_lpi_1_dfm_mx0,
          and_102_nl);
      pixel_processing_if_pixel_processing_if_if_nor_itm_2 <= pixel_processing_if_pixel_processing_if_if_nor_itm;
      system_input_output_vld_sva_dfm_st_2 <= system_input_output_vld_sva_dfm_st_1;
      else_io_read_in_data_vld_rsc_svs_st_2 <= else_io_read_in_data_vld_rsc_svs_st_1;
      asn_itm_1 <= asn_itm;
      main_stage_0_2 <= ~ (fsm_output[2]);
      buffer_slc_buffer_c_5_0_1_itm_2 <= system_input_c_sva[5:0];
      buffer_acc_3_itm_2 <= nl_buffer_acc_3_itm_2[3:0];
      buffer_acc_1_itm_2 <= nl_buffer_acc_1_itm_2[3:0];
      else_io_read_in_data_vld_rsc_svs <= MUX_s_1_2_2(in_data_vld_rsci_d, else_io_read_in_data_vld_rsc_svs,
          or_tmp_56);
      clip_window_switch_lp_3_asn_2_itm <= system_input_window_8_sva;
      system_input_din_sva_1 <= in_data_rsci_d;
      buffer_t0_sva_1 <= buffer_buf_rsci_q_d;
      if_if_if_and_mdf_sva_2 <= if_if_if_and_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      buffer_buf_vinit_ndx_sva <= 10'b1001111111;
    end
    else if ( fsm_output[2] ) begin
      buffer_buf_vinit_ndx_sva <= buffer_buf_acc_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_window_6_sva <= 3'b0;
      system_input_window_7_sva <= 3'b0;
    end
    else if ( or_tmp_42 ) begin
      system_input_window_6_sva <= buffer_qr_lpi_1_dfm_mx0;
      system_input_window_7_sva <= buffer_qr_1_lpi_1_dfm_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_window_8_sva <= 3'b0;
    end
    else if ( and_2_cse & (fsm_output[4]) ) begin
      system_input_window_8_sva <= in_data_rsci_d;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      pixel_processing_threshold_sva <= 3'b100;
    end
    else if ( and_itm & (fsm_output[5]) ) begin
      pixel_processing_threshold_sva <= mcu_data_rsci_q_d[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_r_sva <= 32'b0;
    end
    else if ( ~(or_dcpl | system_input_system_input_nand_tmp | (~ (fsm_output[3])))
        ) begin
      system_input_r_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000, (system_input_if_2_qelse_acc_nl),
          (system_input_if_2_system_input_if_2_nand_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      pixel_processing_frame_sva <= 9'b1;
    end
    else if ( (~ or_dcpl) & system_input_system_input_or_tmp & clip_window_clip_window_and_1_tmp
        & clip_window_clip_window_and_tmp & (fsm_output[3]) ) begin
      pixel_processing_frame_sva <= nl_pixel_processing_frame_sva[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_window_4_sva <= 3'b0;
    end
    else if ( ~ or_tmp_48 ) begin
      system_input_window_4_sva <= system_input_window_7_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_window_3_sva <= 3'b0;
    end
    else if ( ~ or_tmp_48 ) begin
      system_input_window_3_sva <= system_input_window_6_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_window_5_sva <= 3'b0;
    end
    else if ( ~ or_tmp_48 ) begin
      system_input_window_5_sva <= system_input_window_8_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_r_filter_sva <= 32'b0;
    end
    else if ( ~(or_dcpl | (~(system_input_system_input_or_tmp & clip_window_clip_window_and_1_tmp))
        | (~ (fsm_output[3]))) ) begin
      system_input_r_filter_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          (system_input_if_1_qelse_acc_nl), (clip_window_switch_lp_2_not_4_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_c_filter_sva <= 32'b0;
    end
    else if ( ~ or_tmp_48 ) begin
      system_input_c_filter_sva <= system_input_c_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_c_sva <= 32'b0;
    end
    else if ( ~ or_tmp_48 ) begin
      system_input_c_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000, (system_input_else_2_acc_nl),
          system_input_system_input_nand_tmp);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_output_vld_sva <= 1'b0;
    end
    else if ( reg_system_input_system_input_output_vld_and_cse ) begin
      system_input_output_vld_sva <= system_input_system_input_or_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      mcu_ready_sva <= 1'b0;
    end
    else if ( fsm_output[5] ) begin
      mcu_ready_sva <= if_if_if_and_tmp | mcu_ready_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      pixel_processing_if_pixel_processing_if_if_nor_itm <= 1'b0;
      system_input_output_vld_sva_dfm_st_1 <= 1'b0;
      else_io_read_in_data_vld_rsc_svs_st_1 <= 1'b0;
    end
    else if ( reg_pixel_processing_if_pixel_processing_if_if_pixel_processing_if_if_and_cse
        ) begin
      pixel_processing_if_pixel_processing_if_if_nor_itm <= ~((pixel_processing_if_if_acc_tmp!=3'b000)
          | (pixel_processing_frame_sva[0]));
      system_input_output_vld_sva_dfm_st_1 <= system_input_system_input_or_tmp;
      else_io_read_in_data_vld_rsc_svs_st_1 <= in_data_vld_rsci_d;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      pixel_processing_if_asn_itm <= 3'b0;
    end
    else if ( mcu_ready_sva & (fsm_output[5]) ) begin
      pixel_processing_if_asn_itm <= pixel_processing_threshold_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      median_max_7_lpi_1_dfm <= 3'b0;
    end
    else if ( (mcu_ready_sva & L1b_if_acc_15_itm_3 & (fsm_output[5])) | and_104_rgt
        ) begin
      median_max_7_lpi_1_dfm <= MUX_v_3_2_2(median_max2_7_lpi_1_dfm_mx0, median_max2_8_lpi_1_dfm_mx0,
          and_104_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      median_max_5_3_lpi_1_dfm <= 3'b0;
      median_max_6_lpi_1_dfm <= 3'b0;
    end
    else if ( reg_median_median_max_or_2_cse ) begin
      median_max_5_3_lpi_1_dfm <= MUX_v_3_2_2(median_max2_5_3_lpi_1_dfm_mx0, L1b_asn_4_mx1w1,
          median_max_and_7_rgt);
      median_max_6_lpi_1_dfm <= MUX_v_3_2_2(L1b_asn_4_mx1w1, median_max2_5_3_lpi_1_dfm_mx0,
          median_max_and_7_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      median_max_4_1_lpi_1_dfm <= 3'b0;
    end
    else if ( (mcu_ready_sva & L1b_if_acc_13_itm_3 & (fsm_output[5])) | and_108_rgt
        ) begin
      median_max_4_1_lpi_1_dfm <= MUX_v_3_2_2(median_max2_4_lpi_1_dfm_mx0, median_max_2_lpi_1_dfm_mx0,
          and_108_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      buffer_sel_1_0_sva_1 <= 1'b0;
    end
    else if ( reg_system_input_system_input_output_vld_and_cse | (fsm_output[2])
        ) begin
      buffer_sel_1_0_sva_1 <= buffer_sel_1_0_sva_dfm_mx0 | (~(mcu_ready_sva & (fsm_output[3])));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      asn_itm <= 1'b0;
    end
    else if ( (fsm_output[6]) | (fsm_output[2]) ) begin
      asn_itm <= mcu_ready_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      clip_window_last_row_0_sva_7 <= 1'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      clip_window_last_row_0_sva_7 <= clip_window_clip_window_and_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      pixel_processing_if_if_1_asn_itm <= 9'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      pixel_processing_if_if_1_asn_itm <= pixel_processing_frame_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      pixel_processing_if_if_1_pixel_processing_if_if_1_if_and_svs_1 <= 1'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      pixel_processing_if_if_1_pixel_processing_if_if_1_if_and_svs_1 <= pixel_processing_if_if_1_pixel_processing_if_if_1_if_and_svs;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_land_1_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      system_input_land_1_lpi_1_dfm_1 <= system_input_land_1_lpi_1_dfm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      median_max2_1_lpi_1_dfm <= 3'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      median_max2_1_lpi_1_dfm <= MUX_v_3_2_2(median_max2_0_lpi_1_dfm_1_mx0, median_max_1_2_lpi_1_dfm_mx0,
          median_max2_and_5_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      median_max_2_2_lpi_1_dfm <= 3'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      median_max_2_2_lpi_1_dfm <= MUX_v_3_2_2(L1b_asn_44_mx0w1, median_max2_2_2_lpi_1_dfm_mx0,
          median_max_and_3_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      median_max2_3_2_lpi_1_dfm <= 3'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      median_max2_3_2_lpi_1_dfm <= MUX_v_3_2_2(median_max_2_1_lpi_1_dfm_mx0, median_max_3_1_lpi_1_dfm_mx0,
          median_max2_and_3_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      median_max_4_2_lpi_1_dfm <= 3'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      median_max_4_2_lpi_1_dfm <= MUX_v_3_2_2(median_max2_3_1_lpi_1_dfm_mx0, median_max2_4_1_lpi_1_dfm_mx0,
          median_max_and_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      median_max2_5_1_lpi_1_dfm <= 3'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      median_max2_5_1_lpi_1_dfm <= MUX_v_3_2_2(system_input_window_8_sva, system_input_window_7_sva,
          median_max2_median_max2_nor_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      clip_window_first_row_0_sva_5 <= 1'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      clip_window_first_row_0_sva_5 <= clip_window_clip_window_nor_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      clip_window_last_col_0_sva_3 <= 1'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      clip_window_last_col_0_sva_3 <= clip_window_clip_window_and_1_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_output_vld_sva_dfm <= 1'b0;
    end
    else if ( ~ or_tmp_56 ) begin
      system_input_output_vld_sva_dfm <= system_input_system_input_or_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      buffer_sel_1_0_sva_dfm <= 1'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      buffer_sel_1_0_sva_dfm <= buffer_sel_1_0_sva_dfm_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      and_2_cse <= 1'b0;
    end
    else if ( fsm_output[3] ) begin
      and_2_cse <= and_2_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      and_itm <= 1'b0;
    end
    else if ( fsm_output[3] ) begin
      and_itm <= pixel_processing_if_if_1_pixel_processing_if_if_1_if_and_svs & system_input_land_1_lpi_1_dfm
          & system_input_system_input_or_tmp & in_data_vld_rsci_d & mcu_ready_sva;
    end
  end
  assign nl_buffer_buf_acc_itm_2  = buffer_buf_vinit_ndx_sva + 10'b1111111111;
  assign and_102_nl = and_dcpl_11 & (~ z_out_1_3);
  assign nl_buffer_acc_3_itm_2  = conv_u2u_3_4({buffer_sel_1_0_sva_dfm_mx0 , 1'b0
      , buffer_sel_1_0_sva_dfm_mx0}) + (system_input_c_sva[9:6]);
  assign nl_buffer_acc_1_itm_2  = (system_input_c_sva[9:6]) + 4'b101;
  assign nl_system_input_if_2_qelse_acc_nl = system_input_r_sva + 32'b1;
  assign system_input_if_2_qelse_acc_nl = nl_system_input_if_2_qelse_acc_nl[31:0];
  assign system_input_if_2_system_input_if_2_nand_nl = ~((system_input_r_sva==32'b00000000000000000000000011101111));
  assign nl_pixel_processing_frame_sva  = pixel_processing_frame_sva + 9'b1;
  assign nl_system_input_if_1_qelse_acc_nl = system_input_r_filter_sva + 32'b1;
  assign system_input_if_1_qelse_acc_nl = nl_system_input_if_1_qelse_acc_nl[31:0];
  assign clip_window_switch_lp_2_not_4_nl = ~ clip_window_clip_window_and_tmp;
  assign nl_system_input_else_2_acc_nl = system_input_c_sva + 32'b1;
  assign system_input_else_2_acc_nl = nl_system_input_else_2_acc_nl[31:0];
  assign median_max2_and_5_nl = z_out_3 & (~ (fsm_output[4]));
  assign median_max_and_3_nl = z_out_1_3 & (~ (fsm_output[4]));
  assign median_max2_and_3_nl = z_out_5_3 & (~ (fsm_output[4]));
  assign median_max_and_1_nl = z_out_6_3 & (~ (fsm_output[4]));
  assign median_max2_median_max2_nor_nl = ~((~(clip_window_clip_window_and_tmp |
      (~ z_out_2_3))) | (fsm_output[4]));
  assign thresholding_if_mux1h_3_nl = MUX1HOT_v_3_3_2((~ pixel_processing_if_asn_itm),
      median_max2_0_lpi_1_dfm_1_mx0, median_max_8_lpi_1_dfm_mx0, {(fsm_output[6])
      , (fsm_output[3]) , (fsm_output[5])});
  assign thresholding_if_mux1h_4_nl = MUX1HOT_v_3_3_2(median_max_5_lpi_1_dfm_mx0,
      (~ median_max_1_2_lpi_1_dfm_mx0), (~ median_max2_9_lpi_1_dfm_1_mx0), {(fsm_output[6])
      , (fsm_output[3]) , (fsm_output[5])});
  assign nl_acc_nl = ({1'b1 , (thresholding_if_mux1h_3_nl) , 1'b1}) + conv_u2u_4_5({(thresholding_if_mux1h_4_nl)
      , 1'b1});
  assign acc_nl = nl_acc_nl[4:0];
  assign z_out_3 = readslicef_5_1_4((acc_nl));
  assign L1b_if_mux1h_3_nl = MUX1HOT_v_3_3_2(median_max2_1_lpi_1_dfm, median_max2_5_lpi_1_dfm_mx0,
      L1b_asn_44_mx0w1, {(fsm_output[5]) , (fsm_output[6]) , (fsm_output[3])});
  assign L1b_if_mux1h_4_nl = MUX1HOT_v_3_3_2((~ median_max2_2_lpi_1_dfm_mx0), (~
      median_max2_6_lpi_1_dfm_mx0), (~ median_max2_2_2_lpi_1_dfm_mx0), {(fsm_output[5])
      , (fsm_output[6]) , (fsm_output[3])});
  assign nl_acc_1_nl = ({1'b1 , (L1b_if_mux1h_3_nl) , 1'b1}) + conv_u2u_4_5({(L1b_if_mux1h_4_nl)
      , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[4:0];
  assign z_out_1_3 = readslicef_5_1_4((acc_1_nl));
  assign L1a_if_mux1h_6_nl = MUX1HOT_v_3_3_2(median_max_6_lpi_1_dfm, system_input_window_7_sva,
      median_max2_7_1_lpi_1_dfm_mx0, {(fsm_output[6]) , (fsm_output[3]) , (fsm_output[5])});
  assign clip_window_mux_2_nl = MUX_v_3_2_2(system_input_window_8_sva, system_input_window_7_sva,
      clip_window_clip_window_and_tmp);
  assign L1a_if_mux1h_7_nl = MUX1HOT_v_3_3_2((~ median_max_7_lpi_1_dfm), (~ (clip_window_mux_2_nl)),
      (~ pixel_processing_window_8_lpi_1_dfm), {(fsm_output[6]) , (fsm_output[3])
      , (fsm_output[5])});
  assign nl_acc_2_nl = ({1'b1 , (L1a_if_mux1h_6_nl) , 1'b1}) + conv_u2u_4_5({(L1a_if_mux1h_7_nl)
      , 1'b1});
  assign acc_2_nl = nl_acc_2_nl[4:0];
  assign z_out_2_3 = readslicef_5_1_4((acc_2_nl));
  assign L1a_if_mux1h_8_nl = MUX1HOT_v_3_3_2(median_max_4_1_lpi_1_dfm, pixel_processing_window_0_lpi_1_dfm,
      median_max_4_2_lpi_1_dfm, {(fsm_output[6]) , (fsm_output[3]) , (fsm_output[5])});
  assign L1a_if_mux1h_9_nl = MUX1HOT_v_3_3_2((~ median_max_5_3_lpi_1_dfm), (~ clip_window_qr_lpi_1_dfm_mx0),
      (~ median_max_5_2_lpi_1_dfm_mx0), {(fsm_output[6]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_acc_3_nl = ({1'b1 , (L1a_if_mux1h_8_nl) , 1'b1}) + conv_u2u_4_5({(L1a_if_mux1h_9_nl)
      , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[4:0];
  assign z_out_3_3 = readslicef_5_1_4((acc_3_nl));
  assign L1a_if_mux_9_nl = MUX_v_3_2_2(pixel_processing_window_2_lpi_1_dfm, median_max2_5_1_lpi_1_dfm,
      fsm_output[5]);
  assign L1a_if_mux_10_nl = MUX_v_3_2_2((~ clip_window_qr_3_lpi_1_dfm_mx0), (~ median_max2_6_1_lpi_1_dfm_mx0),
      fsm_output[5]);
  assign nl_acc_4_nl = ({1'b1 , (L1a_if_mux_9_nl) , 1'b1}) + conv_u2u_4_5({(L1a_if_mux_10_nl)
      , 1'b1});
  assign acc_4_nl = nl_acc_4_nl[4:0];
  assign z_out_4_3 = readslicef_5_1_4((acc_4_nl));
  assign L1a_if_mux_11_nl = MUX_v_3_2_2(median_max_2_1_lpi_1_dfm_mx0, median_max2_5_2_lpi_1_dfm_mx0,
      fsm_output[5]);
  assign L1a_if_mux_12_nl = MUX_v_3_2_2((~ median_max_3_1_lpi_1_dfm_mx0), (~ median_max_7_1_lpi_1_dfm_mx0),
      fsm_output[5]);
  assign nl_acc_5_nl = ({1'b1 , (L1a_if_mux_11_nl) , 1'b1}) + conv_u2u_4_5({(L1a_if_mux_12_nl)
      , 1'b1});
  assign acc_5_nl = nl_acc_5_nl[4:0];
  assign z_out_5_3 = readslicef_5_1_4((acc_5_nl));
  assign L1b_if_mux_6_nl = MUX_v_3_2_2(median_max2_3_1_lpi_1_dfm_mx0, median_max2_3_2_lpi_1_dfm,
      fsm_output[5]);
  assign L1b_if_mux_7_nl = MUX_v_3_2_2((~ median_max2_4_1_lpi_1_dfm_mx0), (~ median_max2_4_2_lpi_1_dfm_mx0),
      fsm_output[5]);
  assign nl_acc_6_nl = ({1'b1 , (L1b_if_mux_6_nl) , 1'b1}) + conv_u2u_4_5({(L1b_if_mux_7_nl)
      , 1'b1});
  assign acc_6_nl = nl_acc_6_nl[4:0];
  assign z_out_6_3 = readslicef_5_1_4((acc_6_nl));
  assign L1a_if_mux_13_nl = MUX_v_3_2_2(median_max2_0_lpi_1_dfm_mx0, median_max_2_2_lpi_1_dfm,
      fsm_output[5]);
  assign L1a_if_mux_14_nl = MUX_v_3_2_2((~ median_max_1_1_lpi_1_dfm_mx0), (~ median_max_3_lpi_1_dfm_mx0),
      fsm_output[5]);
  assign nl_acc_7_nl = ({1'b1 , (L1a_if_mux_13_nl) , 1'b1}) + conv_u2u_4_5({(L1a_if_mux_14_nl)
      , 1'b1});
  assign acc_7_nl = nl_acc_7_nl[4:0];
  assign z_out_7_3 = readslicef_5_1_4((acc_7_nl));
  assign L1b_if_mux_8_nl = MUX_v_3_2_2(median_max2_1_1_lpi_1_dfm_mx0, median_max_6_2_lpi_1_dfm_mx0,
      fsm_output[5]);
  assign L1b_if_mux_9_nl = MUX_v_3_2_2((~ median_max2_2_1_lpi_1_dfm_mx0), (~ median_max2_8_1_lpi_1_dfm_mx0),
      fsm_output[5]);
  assign nl_acc_8_nl = ({1'b1 , (L1b_if_mux_8_nl) , 1'b1}) + conv_u2u_4_5({(L1b_if_mux_9_nl)
      , 1'b1});
  assign acc_8_nl = nl_acc_8_nl[4:0];
  assign z_out_8_3 = readslicef_5_1_4((acc_8_nl));

  function [31:0] MUX1HOT_v_32_4_2;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [3:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    MUX1HOT_v_32_4_2 = result;
  end
  endfunction


  function [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction


  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function  [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function  [2:0] conv_s2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_s2u_2_3 = {vector[1], vector};
  end
  endfunction


  function  [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction


  function  [2:0] conv_u2u_1_3 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_3 = {{2{1'b0}}, vector};
  end
  endfunction


  function  [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function  [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function  [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction

endmodule
`endif

// ------------------------------------------------------------------
//  Design Unit:    filter
// ------------------------------------------------------------------


`ifdef filter
`else
`define filter
module filter (
  clk, rst, in_data_rsc_z, in_data_rsc_lz, in_data_vld_rsc_z, out_data_rsc_z, out_data_rsc_lz,
      mcu_data_rsc_adr, mcu_data_rsc_q, mcu_data_rsc_d, mcu_data_rsc_we
);
  input clk;
  input rst;
  input [2:0] in_data_rsc_z;
  output in_data_rsc_lz;
  input in_data_vld_rsc_z;
  output [2:0] out_data_rsc_z;
  output out_data_rsc_lz;
  output [8:0] mcu_data_rsc_adr;
  input [31:0] mcu_data_rsc_q;
  output [31:0] mcu_data_rsc_d;
  output mcu_data_rsc_we;


  // Interconnect Declarations
  wire [8:0] mcu_data_rsci_adr_d;
  wire [31:0] mcu_data_rsci_d_d;
  wire mcu_data_rsci_we_d;
  wire [31:0] mcu_data_rsci_q_d;
  wire mcu_data_rsci_ram_rw_A_internal_RMASK_B_d;
  wire [9:0] buffer_buf_rsci_radr_d;
  wire [9:0] buffer_buf_rsci_wadr_d;
  wire [2:0] buffer_buf_rsci_d_d;
  wire buffer_buf_rsci_we_d;
  wire buffer_buf_rsci_re_d;
  wire [2:0] buffer_buf_rsci_q_d;
  wire buffer_buf_rsc_we;
  wire [2:0] buffer_buf_rsc_d;
  wire [9:0] buffer_buf_rsc_wadr;
  wire buffer_buf_rsc_re;
  wire [2:0] buffer_buf_rsc_q;
  wire [9:0] buffer_buf_rsc_radr;


  // Interconnect Declarations for Component Instantiations 
  BLOCK_1R1W_RBW #(.data_width(32'sd3),
  .addr_width(32'sd10),
  .depth(32'sd640)) buffer_buf_rsc_comp (
      .radr(buffer_buf_rsc_radr),
      .wadr(buffer_buf_rsc_wadr),
      .d(buffer_buf_rsc_d),
      .we(buffer_buf_rsc_we),
      .re(buffer_buf_rsc_re),
      .clk(clk),
      .q(buffer_buf_rsc_q)
    );
  Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_32_9_512_4_gen mcu_data_rsci (
      .we(mcu_data_rsc_we),
      .d(mcu_data_rsc_d),
      .q(mcu_data_rsc_q),
      .adr(mcu_data_rsc_adr),
      .adr_d(mcu_data_rsci_adr_d),
      .d_d(mcu_data_rsci_d_d),
      .we_d(mcu_data_rsci_we_d),
      .q_d(mcu_data_rsci_q_d),
      .ram_rw_A_internal_RMASK_B_d(mcu_data_rsci_ram_rw_A_internal_RMASK_B_d)
    );
  Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_3_10_640_7_gen buffer_buf_rsci (
      .we(buffer_buf_rsc_we),
      .d(buffer_buf_rsc_d),
      .wadr(buffer_buf_rsc_wadr),
      .re(buffer_buf_rsc_re),
      .q(buffer_buf_rsc_q),
      .radr(buffer_buf_rsc_radr),
      .radr_d(buffer_buf_rsci_radr_d),
      .wadr_d(buffer_buf_rsci_wadr_d),
      .d_d(buffer_buf_rsci_d_d),
      .we_d(buffer_buf_rsci_we_d),
      .re_d(buffer_buf_rsci_re_d),
      .q_d(buffer_buf_rsci_q_d)
    );
  filter_core filter_core_inst (
      .clk(clk),
      .rst(rst),
      .in_data_rsc_z(in_data_rsc_z),
      .in_data_rsc_lz(in_data_rsc_lz),
      .in_data_vld_rsc_z(in_data_vld_rsc_z),
      .out_data_rsc_z(out_data_rsc_z),
      .out_data_rsc_lz(out_data_rsc_lz),
      .mcu_data_rsci_adr_d(mcu_data_rsci_adr_d),
      .mcu_data_rsci_d_d(mcu_data_rsci_d_d),
      .mcu_data_rsci_we_d(mcu_data_rsci_we_d),
      .mcu_data_rsci_q_d(mcu_data_rsci_q_d),
      .mcu_data_rsci_ram_rw_A_internal_RMASK_B_d(mcu_data_rsci_ram_rw_A_internal_RMASK_B_d),
      .buffer_buf_rsci_radr_d(buffer_buf_rsci_radr_d),
      .buffer_buf_rsci_wadr_d(buffer_buf_rsci_wadr_d),
      .buffer_buf_rsci_d_d(buffer_buf_rsci_d_d),
      .buffer_buf_rsci_we_d(buffer_buf_rsci_we_d),
      .buffer_buf_rsci_re_d(buffer_buf_rsci_re_d),
      .buffer_buf_rsci_q_d(buffer_buf_rsci_q_d)
    );
endmodule
`endif



