
//------> C:/PROGRA~1/MENTOR~1/CATAPU~1.0C/Mgc_home/pkgs/siflibs/mgc_in_wire_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


`ifdef mgc_in_wire_v1
`else
`define mgc_in_wire_v1
module mgc_in_wire_v1 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] d;
  input  [width-1:0] z;

  wire   [width-1:0] d;

  assign d = z;

endmodule
`endif


//------> C:/PROGRA~1/MENTOR~1/CATAPU~1.0C/Mgc_home/pkgs/siflibs/mgc_out_stdreg_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

`ifdef mgc_out_stdreg_v1
`else
`define mgc_out_stdreg_v1
module mgc_out_stdreg_v1 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule
`endif




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0c/745553 Production Release
//  HLS Date:       Wed Oct 11 16:38:17 PDT 2017
// 
//  Generated by:   Fitkit@DESKTOP-NJUNEBJ
//  Generated date: Tue Oct 31 12:27:20 2017
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    genpix_core
// ------------------------------------------------------------------


`ifdef genpix_core
`else
`define genpix_core
module genpix_core (
  clk, rst, pause_rsc_z, req_rsc_z, pixel_rsc_z, pixel_vld_rsc_z
);
  input clk;
  input rst;
  input pause_rsc_z;
  input req_rsc_z;
  output [2:0] pixel_rsc_z;
  output pixel_vld_rsc_z;


  // Interconnect Declarations
  wire pause_rsci_d;
  wire req_rsci_d;
  reg [2:0] pixel_rsci_d;
  reg pixel_vld_rsci_d;
  wire not_tmp_14;
  wire or_dcpl_16;
  wire or_dcpl_17;
  reg [8:0] r_sva;
  reg [8:0] c_sva;
  reg [8:0] base_r_sva;
  wire [9:0] nl_base_r_sva;
  reg [8:0] base_c_sva;
  wire [9:0] nl_base_c_sva;
  reg [9:0] noise_cnt_sva;
  reg [5:0] frame_cnt_sva;
  wire [6:0] nl_frame_cnt_sva;
  reg update_base_pos_inc_r_1_sva;
  reg update_base_pos_inc_c_1_sva;
  reg if_1_asn_itm;
  wire [8:0] diff_c_sva;
  wire [9:0] nl_diff_c_sva;
  wire [8:0] diff_r_sva;
  wire [9:0] nl_diff_r_sva;
  wire [3:0] diff_aux_sva;
  wire [4:0] nl_diff_aux_sva;
  wire reg_update_base_pos_update_base_pos_inc_c_nor_cse;
  wire if_acc_tmp_3;
  wire equal_cse_sva;
  wire if_1_if_unequal_tmp;
  wire if_1_unequal_tmp;
  wire update_base_pos_inc_c_1_sva_dfm;
  wire update_base_pos_inc_r_1_sva_dfm;
  wire aelse_acc_itm_3;

  wire[3:0] aelse_acc_nl;
  wire[4:0] nl_aelse_acc_nl;
  wire[3:0] if_acc_nl;
  wire[4:0] nl_if_acc_nl;
  wire[2:0] and_1_nl;
  wire[0:0] if_if_and_nl;
  wire[0:0] or_20_nl;
  wire[8:0] if_1_if_else_acc_nl;
  wire[9:0] nl_if_1_if_else_acc_nl;
  wire[8:0] if_1_else_acc_nl;
  wire[9:0] nl_if_1_else_acc_nl;
  wire[9:0] if_1_qelse_acc_nl;
  wire[10:0] nl_if_1_qelse_acc_nl;
  wire[0:0] not_5_nl;
  wire[2:0] mux_nl;
  wire[9:0] acc_7_nl;
  wire[11:0] nl_acc_7_nl;

  // Interconnect Declarations for Component Instantiations 
  mgc_in_wire_v1 #(.rscid(32'sd1),
  .width(32'sd1)) pause_rsci (
      .d(pause_rsci_d),
      .z(pause_rsc_z)
    );
  mgc_in_wire_v1 #(.rscid(32'sd2),
  .width(32'sd1)) req_rsci (
      .d(req_rsci_d),
      .z(req_rsc_z)
    );
  mgc_out_stdreg_v1 #(.rscid(32'sd3),
  .width(32'sd3)) pixel_rsci (
      .d(pixel_rsci_d),
      .z(pixel_rsc_z)
    );
  mgc_out_stdreg_v1 #(.rscid(32'sd4),
  .width(32'sd1)) pixel_vld_rsci (
      .d(pixel_vld_rsci_d),
      .z(pixel_vld_rsc_z)
    );
  assign nl_aelse_acc_nl = conv_u2u_3_4(diff_r_sva[8:6]) + 4'b1111;
  assign aelse_acc_nl = nl_aelse_acc_nl[3:0];
  assign aelse_acc_itm_3 = readslicef_4_1_3((aelse_acc_nl));
  assign nl_if_acc_nl = conv_u2u_3_4(diff_c_sva[8:6]) + 4'b1111;
  assign if_acc_nl = nl_if_acc_nl[3:0];
  assign if_acc_tmp_3 = readslicef_4_1_3((if_acc_nl));
  assign reg_update_base_pos_update_base_pos_inc_c_nor_cse = ~(if_1_if_unequal_tmp
      | if_1_unequal_tmp | not_tmp_14);
  assign nl_acc_7_nl = ({1'b1 , diff_c_sva}) + conv_u2u_9_10(~ diff_r_sva) + 10'b1;
  assign acc_7_nl = nl_acc_7_nl[9:0];
  assign mux_nl = MUX_v_3_2_2((diff_c_sva[5:3]), (diff_r_sva[5:3]), readslicef_10_1_9((acc_7_nl)));
  assign nl_diff_aux_sva = conv_u2u_3_4(~ (mux_nl)) + conv_u2u_3_4(frame_cnt_sva[5:3]);
  assign diff_aux_sva = nl_diff_aux_sva[3:0];
  assign nl_diff_c_sva = c_sva - base_c_sva;
  assign diff_c_sva = nl_diff_c_sva[8:0];
  assign nl_diff_r_sva = r_sva - base_r_sva;
  assign diff_r_sva = nl_diff_r_sva[8:0];
  assign equal_cse_sva = (noise_cnt_sva==10'b1111110000);
  assign if_1_if_unequal_tmp = ~((r_sva==9'b011101111));
  assign if_1_unequal_tmp = ~((c_sva==9'b100111111));
  assign update_base_pos_inc_c_1_sva_dfm = (update_base_pos_inc_c_1_sva & ((base_c_sva!=9'b000000000)))
      | ((base_c_sva==9'b100000000));
  assign update_base_pos_inc_r_1_sva_dfm = (update_base_pos_inc_r_1_sva & ((base_r_sva!=9'b000000000)))
      | ((base_r_sva==9'b010110000));
  assign not_tmp_14 = ~(if_1_asn_itm | req_rsci_d);
  assign or_dcpl_16 = not_tmp_14 | (c_sva!=9'b100111111);
  assign or_dcpl_17 = or_dcpl_16 | (r_sva!=9'b011101111);
  always @(posedge clk) begin
    if ( rst ) begin
      frame_cnt_sva <= 6'b0;
    end
    else if ( ~ or_dcpl_17 ) begin
      frame_cnt_sva <= nl_frame_cnt_sva[5:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      pixel_rsci_d <= 3'b0;
    end
    else if ( ~ not_tmp_14 ) begin
      pixel_rsci_d <= MUX_v_3_2_2((and_1_nl), 3'b111, (or_20_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      r_sva <= 9'b0;
    end
    else if ( ~ or_dcpl_16 ) begin
      r_sva <= MUX_v_9_2_2(9'b000000000, (if_1_if_else_acc_nl), if_1_if_unequal_tmp);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      c_sva <= 9'b0;
    end
    else if ( ~ not_tmp_14 ) begin
      c_sva <= MUX_v_9_2_2(9'b000000000, (if_1_else_acc_nl), if_1_unequal_tmp);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      noise_cnt_sva <= 10'b0;
    end
    else if ( ~ not_tmp_14 ) begin
      noise_cnt_sva <= MUX_v_10_2_2(10'b0000000000, (if_1_qelse_acc_nl), (not_5_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      pixel_vld_rsci_d <= 1'b0;
      if_1_asn_itm <= 1'b1;
    end
    else begin
      pixel_vld_rsci_d <= ~ pause_rsci_d;
      if_1_asn_itm <= 1'b0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      base_c_sva <= 9'b1100100;
    end
    else if ( ~ or_dcpl_17 ) begin
      base_c_sva <= nl_base_c_sva[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      base_r_sva <= 9'b1100100;
    end
    else if ( ~ or_dcpl_17 ) begin
      base_r_sva <= nl_base_r_sva[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      update_base_pos_inc_c_1_sva <= 1'b0;
      update_base_pos_inc_r_1_sva <= 1'b0;
    end
    else if ( reg_update_base_pos_update_base_pos_inc_c_nor_cse ) begin
      update_base_pos_inc_c_1_sva <= update_base_pos_inc_c_1_sva_dfm;
      update_base_pos_inc_r_1_sva <= update_base_pos_inc_r_1_sva_dfm;
    end
  end
  assign nl_frame_cnt_sva  = frame_cnt_sva + 6'b1;
  assign if_if_and_nl = aelse_acc_itm_3 & if_acc_tmp_3;
  assign and_1_nl = MUX_v_3_2_2(3'b000, (diff_aux_sva[2:0]), (if_if_and_nl));
  assign or_20_nl = (if_acc_tmp_3 & aelse_acc_itm_3 & (diff_aux_sva[3])) | equal_cse_sva;
  assign nl_if_1_if_else_acc_nl = r_sva + 9'b1;
  assign if_1_if_else_acc_nl = nl_if_1_if_else_acc_nl[8:0];
  assign nl_if_1_else_acc_nl = c_sva + 9'b1;
  assign if_1_else_acc_nl = nl_if_1_else_acc_nl[8:0];
  assign nl_if_1_qelse_acc_nl = noise_cnt_sva + 10'b1;
  assign if_1_qelse_acc_nl = nl_if_1_qelse_acc_nl[9:0];
  assign not_5_nl = ~ equal_cse_sva;
  assign nl_base_c_sva  = base_c_sva + conv_s2u_2_9({update_base_pos_inc_c_1_sva_dfm
      , 1'b1});
  assign nl_base_r_sva  = base_r_sva + conv_s2u_2_9({update_base_pos_inc_r_1_sva_dfm
      , 1'b1});

  function [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction


  function  [8:0] conv_s2u_2_9 ;
    input [1:0]  vector ;
  begin
    conv_s2u_2_9 = {{7{vector[1]}}, vector};
  end
  endfunction


  function  [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function  [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction

endmodule
`endif

// ------------------------------------------------------------------
//  Design Unit:    genpix
// ------------------------------------------------------------------


`ifdef genpix
`else
`define genpix
module genpix (
  clk, rst, pause_rsc_z, req_rsc_z, pixel_rsc_z, pixel_vld_rsc_z
);
  input clk;
  input rst;
  input pause_rsc_z;
  input req_rsc_z;
  output [2:0] pixel_rsc_z;
  output pixel_vld_rsc_z;



  // Interconnect Declarations for Component Instantiations 
  genpix_core genpix_core_inst (
      .clk(clk),
      .rst(rst),
      .pause_rsc_z(pause_rsc_z),
      .req_rsc_z(req_rsc_z),
      .pixel_rsc_z(pixel_rsc_z),
      .pixel_vld_rsc_z(pixel_vld_rsc_z)
    );
endmodule
`endif



